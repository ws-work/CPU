`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 2017/11/02 15:12:22
// Design Name:
// Module Name: datapath
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module datapath(input wire clk,rst,
                output wire[31:0] pcF,
                input wire[31:0] instrF,
                input wire pcsrcD,branchD,
                input wire jumpD,
                output wire equalD,
                output wire[5:0] opD,functD,
                input wire memtoregE,
                input wire alusrcE,regdstE,
                input wire regwriteE,
                input wire[5:0] alucontrolE,
                output wire flushE,
                input wire memtoregM,
                input wire regwriteM,
                output wire[31:0] aluoutM,writedataM,
                input wire[31:0] readdataM,
                input wire memtoregW,
                input wire regwriteW);

    //fetch stage
    wire stallF;
    //FD
    wire [31:0] pcnextFD,pcnextbrFD,pcplus4F,pcbranchD;
    //decode stage
    wire [31:0] pcplus4D,instrD;
    wire forwardaD,forwardbD;
    wire [4:0] rsD,rtD,rdD,saD;
    wire flushD,stallD;
    wire [31:0] signimmD,signimmshD;
    wire [31:0] srcaD,srca2D,srcbD,srcb2D;
    //execute stage
    wire [1:0] forwardaE,forwardbE;
    wire [4:0] rsE,rtE,rdE,saE;
    wire [4:0] writeregE;
    wire [31:0] signimmE;
    wire [31:0] srcaE,srca2E,srcbE,srcb2E,srcb3E;
    wire [31:0] aluoutE;
    //mem stage
    wire [4:0] writeregM;
    //writeback stage
    wire [4:0] writeregW;
    wire [31:0] aluoutW,readdataW,resultW;
    wire divstallE;
    wire overflowE,zeroE;
    wire [63:0] aluoutE_64;
    wire [31:0] hi_o;
    wire [31:0] lo_o;
    wire hilo_ena;

    //hazard detection
    hazard h(
    //fetch stage
    stallF,
    //decode stage
    rsD,rtD,
    branchD,
    forwardaD,forwardbD,
    stallD,
    //execute stage
    rsE,rtE,
    writeregE,
    regwriteE,
    memtoregE,
    forwardaE,forwardbE,
    flushE,
    //mem stage
    writeregM,
    regwriteM,
    memtoregM,
    //write back stage
    writeregW,
    regwriteW
    );

    //next PC logic (operates in fetch an decode)
    mux2 #(32) pcbrmux(pcplus4F,pcbranchD,pcsrcD,pcnextbrFD);
    mux2 #(32) pcmux(pcnextbrFD,
    {pcplus4D[31:28],instrD[25:0],2'b00},
    jumpD,pcnextFD);

    //regfile (operates in decode and writeback)
    regfile rf(clk,regwriteW,rsD,rtD,writeregW,resultW,srcaD,srcbD);

    //fetch stage logic
    pc #(32) pcreg(clk,rst,~stallF,pcnextFD,pcF);
    adder pcadd1(pcF,32'b100,pcplus4F);
    //decode stage
    flopenr #(32) r1D(clk,rst,~stallD,pcplus4F,pcplus4D);
    flopenrc #(32) r2D(clk,rst,~stallD,flushD,instrF,instrD);
    signext se(instrD[15:0],signimmD);
    sl2 immsh(signimmD,signimmshD);
    adder pcadd2(pcplus4D,signimmshD,pcbranchD);
    mux2 #(32) forwardamux(srcaD,aluoutM,forwardaD,srca2D);
    mux2 #(32) forwardbmux(srcbD,aluoutM,forwardbD,srcb2D);
    eqcmp comp(srca2D,srcb2D,equalD);

    assign opD    = instrD[31:26];
    assign functD = instrD[5:0];
    assign rsD    = instrD[25:21];
    assign rtD    = instrD[20:16];
    assign rdD    = instrD[15:11];
    assign saD    = instrD[10:6];

    //execute stage
    floprc #(32) r1E(clk,rst,flushE,srcaD,srcaE);
    floprc #(32) r2E(clk,rst,flushE,srcbD,srcbE);
    floprc #(32) r3E(clk,rst,flushE,signimmD,signimmE);
    floprc #(5) r4E(clk,rst,flushE,rsD,rsE);
    floprc #(5) r5E(clk,rst,flushE,rtD,rtE);
    floprc #(5) r6E(clk,rst,flushE,rdD,rdE);
    floprc #(5) r7E(clk,rst,flushE,saD,saE);

    mux3 #(32) forwardaemux(srcaE,resultW,aluoutM,forwardaE,srca2E);
    mux3 #(32) forwardbemux(srcbE,resultW,aluoutM,forwardbE,srcb2E);
    mux2 #(32) srcbmux(srcb2E,signimmE,alusrcE,srcb3E);//b��1��imm��reg
    //div div(clk,rsk,0,);
    alu alu(
    .a(srca2E),
    .b(srcb3E),
    .sa(saE),
    .op(alucontrolE),
    .lo_o(lo_o),
    .hi_o(hi_o),
    .y(aluoutE),
    .overflow(overflowE),
    .zero(zeroE),
    .hilo_ena(hilo_ena),
    .hilo(aluoutE_64)
    );

    hilo_reg hilo_reg(
        .clk(clk),
        .rst(rst),
        .we(hilo_ena),
        .hi_i(aluoutE_64[63:32]),
        .lo_i(aluoutE_64[31:0]),
        .hi_o(hi_o),
        .lo_o(lo_o)
    );

    mux2 #(5) wrmux(rtE,rdE,regdstE,writeregE);

    //mem stage
    flopr #(32) r1M(clk,rst,srcb2E,writedataM);
    flopr #(32) r2M(clk,rst,aluoutE,aluoutM);
    flopr #(5) r3M(clk,rst,writeregE,writeregM);

    //writeback stage
    flopr #(32) r1W(clk,rst,aluoutM,aluoutW);
    flopr #(32) r2W(clk,rst,readdataM,readdataW);
    flopr #(5) r3W(clk,rst,writeregM,writeregW);
    mux2 #(32) resmux(aluoutW,readdataW,memtoregW,resultW);
endmodule
